/* Name: Mohammed Abdul Haq
UVM Test-Bench Name: AHBLite_APB_Bridge
*/
`include "sequence_item_0.sv"
`include "sequence_0.sv"
`include "sequencer_0.sv"
`include "driver_0.sv"
`include "monitor_0.sv"
`include "agent_0.sv"

`include "sequence_item_1.sv"
`include "sequence_1.sv"
`include "sequencer_1.sv"
`include "driver_1.sv"
`include "monitor_1.sv"
`include "agent_1.sv"

`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"
